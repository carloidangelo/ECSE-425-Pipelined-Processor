--Instruction_Memory.vhd