--PipelinedProcessor.vhd