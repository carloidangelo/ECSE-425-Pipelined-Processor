--Fetch.vhd