-- OPCODE signal for ALU operations 

--    R-Type
-- add = "00000";
-- and = "00001";
-- div = "00010";
-- nor = "00011";
-- or = "00100";
-- slt = "00101";
-- sub = "00110";
-- xor = "00111";
-- mult = "01000";      
-- mfhi = "01001";
-- mflo = "01010";
-- sra = "01011";
-- sll = "01100";
-- srl = "01101";
-- jr = "01110";
 
--    Jtype
-- j = "01111";
-- jal = "10000";       

--     Itype
-- addi = "10001";
-- andi = "10010";
-- ori = "10011";
-- xori = "10100";
-- lw = "10101";
-- lui = "10110";
-- sw = "10111";
-- slti = "11000";
-- beq = "11001";
-- bne = "11010";
