--Execute.vhd