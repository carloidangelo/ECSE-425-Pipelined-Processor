--Write_Back.vhd