--Decode.vhd