--Memory.vhd